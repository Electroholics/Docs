** Darlington boost op-amp (from EDN May 29, 1986 pg 133 -> with minor changes)

vin 1 0 sin(0 5 10k) dc 0 ac 1
vcc     11      0       15.0
vee     12      0       -15.0
r1      0       2       10k
r2      2     out       10k
r3      5       6       2k
r4      5      20       33k
r5     20      10       2k
r6     11       7       1.2k
r7     18      12       1.2k
r8     14      15       1k
r9     16      17       1k
r10    15     out       .1
r11    17     out       .1
r12     1       3       5k
rload out       0       8
c1      2       4       39pf
d1     11       6          D1N4148
d2      8       9          D1N4148
d3      9       4          D1N4148
d4      4      13          d1n4148
d5     13      19          d1n4148
d6     10      12          d1n4148
q1      8       5      7   q2n3906
q2     19      20     18   q2n3904
q3      8      14    out   q2n2222A
q4     19      16    out   q2n2907A
x1      3       2     11     12   4  lf156
x2     11       8     15   q2n6384
x3     12      19     17   q2n6649
.include lf156

* Note: this next line are meaningful only in batch mode
.save 1 out
* Note: these next lines are meaningful only in batch mode
* or when the "run" command is given in interactive mode
.AC dec 15 1 100meghz
.tran .5us 200us
.four 10k out
***************************
*  models and subcircuits *
***************************
.MODEL D1N4148 D (IS=14.2P RS=4.2 N=1.7 BV=74.9 IBV=10U
+ CJO=1.73P VJ=.75 M=.333 TT=5.76N)
*   75 Volt  .01 Amp  .004 us  Si Diode  07-08-1991
**********
.MODEL Q2N3906 PNP (IS=8.012404E-17 NF=1 BF=136 VAF=113 IKF=65M
+ ISE=800F NE=2 BR=4 NR=1 VAR=20 IKR=97.5M RE=3.63 RB=14.5
+ RC=1.45 XTB=1.5 CJE=11.8P CJC=8.81P TF=636P TR=95.6N)
*   40 Volt  .2 Amp  250 MHz  SiPNP  Transistor  06-28-1991
**********
.MODEL Q2N3904 NPN (IS=4.667347E-17 NF=1 BF=238 VAF=113 IKF=65M
+ ISE=1.18P NE=2 BR=4 NR=1 VAR=24 IKR=97.5M RE=2.63 RB=10.5
+ RC=1.05 XTB=1.5 CJE=9.46P CJC=7.83P TF=530P TR=85N)
*   40 Volt  .2 Amp  300 MHz  SiNPN  Transistor  06-28-1991
**********
.MODEL Q2N2222A NPN (IS=5.632971E-19 NF=1 BF=175 VAF=113 IKF=.4
+ ISE=237F NE=2 BR=4 NR=1 VAR=24 IKR=.6 RE=.963 RB=3.85
+ RC=.385 XTB=1.5 CJE=29.5P CJC=19.2P TF=530P TR=95.6N)
*   40 Volt  .8 Amp  300 MHz  SiNPN  Transistor  06-28-1991
**********
.MODEL Q2N2907A PNP (IS=1.536728E-18 NF=1 BF=103 VAF=139 IKF=.5
+ ISE=96.0F NE=2 BR=4 NR=1 VAR=20 IKR=.75 RE=1.56 RB=6.25
+ RC=.625 XTB=1.5 CJE=46.0P CJC=19.2P TF=794P TR=34N)
*   60 Volt  .6 Amp  200 MHz  SiPNP  Transistor  06-28-1991
**********
.SUBCKT Q2N6384  1 2 3
*    TERMINALS:  C B E
Q1 1 2 4 QPWR .1
Q2 1 4 3 QPWR
R1 2 4  4K
R2 4 3  50
D1 3 1  DSUB
.MODEL QPWR NPN (IS=12P NF=1 BF=49.3 VAF=139 IKF=7.5
+ ISE=21.2P NE=2 BR=4 NR=1 VAR=20 IKR=11.2 RE=.115 RB=.46
+ RC=46M XTB=1.5 CJE=2.21N CJC=481P TF=1.34P TR=3.67U)
.MODEL DSUB D (IS=12P N=1 RS=.115 BV=60 IBV=.001
+ CJO=481P TT=3.67U)
.ENDS
*   60 Volt  10 Amp  NPN Darlington Transistor  06-28-1991
**********
.SUBCKT Q2N6649  1 2 3
*    TERMINALS:  C B E
Q1 1 2 4 QPWR .1
Q2 1 4 3 QPWR
R1 2 4  4K
R2 4 3  50
D1 1 3  DSUB
.MODEL QPWR PNP (IS=12P NF=1 BF=49.3 VAF=139 IKF=7.5
+ ISE=21.2P NE=2 BR=4 NR=1 VAR=20 IKR=11.2 RE=.115 RB=.46
+ RC=46M XTB=1.5 CJE=2.21N CJC=481P TF=1.34P TR=3.67U)
.MODEL DSUB D (IS=12P N=1 RS=.115 BV=60 IBV=.001
+ CJO=481P TT=3.67U)
.ENDS
*   60 Volt  10 Amp  PNP Darlington Transistor  06-28-1991
.end
